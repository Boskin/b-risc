`include "opcodes.vh"

module tb_instruction_memory;

endmodule
