`ifndef CONFIG_VH
`define CONFIG_VH

`define ADDR_W 32
`define WORD_W 32
`define INSTR_W 32
`define REG_COUNT 32

`endif
