`ifndef MEM_CODES_VH
`define MEM_CODES_VH

`define MEM_COUNT_W

`define MEM_COUNT_NONE 0
`define MEM_COUNT_BYTE 1
`define MEM_COUNT_HALF 2
`define MEM_COUNT_WORD 3

`define MEM_CODE_W 2

`define MEM_CODE_INVALID 0
`define MEM_CODE_READ 1
`define MEM_CODE_WRITE 2
`define MEM_CODE_MISALIGNED 2

`endif
