module id(
    instr,
    
    alu_op,
    
);

endmodule
