`ifndef ALU_OP_VH
`define ALU_OP_VH

// ALU operations
`define ALU_ADD 0
`define ALU_AND 1
`define ALU_OR 2
`define ALU_XOR 3
`define ALU_SLT 4
`define ALU_SLTU 5
`define ALU_SUB 6
`define ALU_SLL 7
`define ALU_SRL 8
`define ALU_SRA 9

`define ALU_OP_W 4

`endif
